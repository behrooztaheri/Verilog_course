module Adder_(
    input [3:0] X,
    input [3:0] Y,
    output [4:0] Z
);

    assign Z = X + Y;

endmodule