module xor_gate(input a, input b, output Out);

    assign Out = a ^ b;

endmodule